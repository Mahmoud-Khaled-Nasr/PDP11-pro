LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE.ALL;

ENTITY GENERAL_REGISTER IS
	GENERIC (SIZE : INTEGER := 32);
	PORT (
		D,DX		: IN STD_LOGIC_VECTOR (SIZE-1 DOWNTO 0);	--DX : IF ENB=1 INPUT=D , IF ENBX=1 INPUT=DX
		CLK,RST,ENB,ENBX: IN STD_LOGIC;
		Q,QX 		: OUT STD_LOGIC_VECTOR (SIZE-1 DOWNTO 0)	--QX IS THE SAME AS 'Q' NO THING ELSE
	);

END ENTITY GENERAL_REGISTER;



architecture GENERAL_REGISTER_ARCH of GENERAL_REGISTER is

SIGNAL SEL :STD_LOGIC;
begin

SEL <= ENB XOR ENBX;

	process(RST,CLK,ENB,ENBX)
	begin
		if (RST='1') then
			Q  <= (OTHERS=>'0');
			QX <= (OTHERS=>'0');
		--Changed from rising edge to falling edge
	elsif(falling_edge(CLK) AND SEL='1')then
			IF(ENB='1') THEN
				Q  <= D;
				QX <= D;
			ELSIF(ENBX='1')THEN
				Q  <= DX;
				QX <= DX;
			END IF;	
		end if;
	end process;


end GENERAL_REGISTER_ARCH;
