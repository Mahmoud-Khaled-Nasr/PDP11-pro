LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE.ALL;

--TODO WHICH BUS USES THE MAR
ENTITY MAR_REGISTER IS
	GENERIC (SIZE : INTEGER := 32);
	PORT (
		DATA_IN_B, DATA_IN_Z : IN STD_LOGIC_VECTOR (SIZE-1 DOWNTO 0);
		CLK : IN STD_LOGIC;
		BUS_B_IN_ENABLE, BUS_B_OUT_ENABLE, BUS_Z_IN_ENABLE : IN STD_LOGIC ;
		DATA_OUT_B : OUT STD_LOGIC_VECTOR (SIZE-1 DOWNTO 0)
	);

END ENTITY MAR_REGISTER;
