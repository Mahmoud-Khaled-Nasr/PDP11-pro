LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE;

ENTITY RAM IS
	GENERIC (ADDRESS_SIZE : INTEGER :=11; CELL_SIZE : INTEGER := 16);	--11BIT FOR MEMORY ADDRESS_SIZE PROVIDES 2K BIT MEMORY
	PORT (
		DATA_IN 	:IN STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
		--TYP : READING MODE 16 BIT IF 0 32 IF 1
		RD, WRT,TYP 	: IN STD_LOGIC;
		CLK,ENB		:IN STD_LOGIC;
		ADDRESS		:IN STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0);
		DATA_OUT 	: OUT STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
		--MDR_READ IS THE SIGNAL TO ENABLE THE MDR TO READ FROM THE MEMORY
		
		MFC, MDR_READ 	:OUT STD_LOGIC
		
	);
END ENTITY RAM;
		

ARCHITECTURE RAM_ARCH OF RAM IS

	TYPE ram_type IS ARRAY(0 TO 2047) OF std_logic_vector(CELL_SIZE-1 DOWNTO 0);
	SIGNAL ram : ram_type ;
	
	BEGIN
		PROCESS(CLK) IS
			BEGIN
				IF rising_edge(clk) THEN  
					IF WRT = '1' THEN
						ram(to_integer(unsigned(ADDRESS))) <= DATA_IN;
					END IF;
				END IF;
		END PROCESS;
		DATA_OUT <= ram(to_integer(unsigned(ADDRESS)));
END RAM_ARCH;