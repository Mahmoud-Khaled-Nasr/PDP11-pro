LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE.ALL;

ENTITY SRC_FETCHING_BLOCK IS
	PORT (
		IR : IN std_logic_vector (IR_SIZE-1 DOWNTO 0);
		INSTRUCTION_COUNTER : IN STD_LOGIC_VECTOR (INSTRUCTION_COUNTER_OUTPUT_SIZE-1 DOWNTO 0); 
		CONTROL_WORD: OUT STD_LOGIC_VECTOR (ROM_WIDTH-1 DOWNTO 0);
		INITIAL_ADDRESS: OUT STD_LOGIC_VECTOR (INSTRUCTION_COUNTER_OUTPUT_SIZE-1 DOWNTO 0) );
END ENTITY SRC_FETCHING_BLOCK;

ARCHITECTURE FETCH_SOURCE OF SRC_FETCHING_BLOCK IS
	-----------------Signals---------
	SIGNAL ROM_OUTPUT : STD_LOGIC_VECTOR(ROM_WIDTH-1 DOWNTO 0);
	SIGNAL IR_SRC : STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL IR_SRC_ADDRESS_MODE : STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL INITIAL_ADDRESS_SIGNAL : STD_LOGIC_VECTOR (INSTRUCTION_COUNTER_OUTPUT_SIZE-1 DOWNTO 0) := "000";
	-----------------ROM------------
	CONSTANT ROM_LENGTH : INTEGER := 8; --LENGTH OF THE ROM USED IN THIS BLOCK
	TYPE ROM_TYPE IS ARRAY(0 TO ROM_LENGTH - 1) OF std_logic_vector(ROM_WIDTH-1 DOWNTO 0);
	CONSTANT ROM_DATA : ROM_TYPE := 
	(
		0 => B"01101_1111_0000_1001_1111_00_10100",
		1 => B"00000_1010_0000_1100_0000_00_00010",
		2 => B"01111_1111_0000_0000_1111_01_10100",
		3 => B"00000_1010_0000_1100_0000_00_00010",
		4 => B"01100_1000_0000_1001_1000_00_10000",
		5 => B"00001_1010_1111_0000_0000_01_10100",
		6 => B"00000_1010_0000_1100_0000_00_00010",
		7 => "ZZZZZZZZZZZZZZZZZZZZZZZZZZZZ"
	);
	BEGIN
	-------------------------Circuit that calculate the initial value-----------
	IR_SRC_ADDRESS_MODE <= IR(11 DOWNTO 9);
	INITIAL_ADDRESS <= "000" WHEN IR_SRC_ADDRESS_MODE = AUTO_INCR_ADDRESSING_MODE 
		ELSE "010" WHEN IR_SRC_ADDRESS_MODE = AUTO_DECR_ADDRESSING_MODE
		ELSE "100" WHEN IR_SRC_ADDRESS_MODE = INDEXED_ADDRESSING_MODE
		ELSE "111";
	-------------------------the ROM process---------------
	ROM_OUTPUT <= ROM_DATA(to_integer(unsigned(INSTRUCTION_COUNTER))) WHEN INSTRUCTION_COUNTER < 8
		ELSE ROM_DATA(to_integer(unsigned(INITIAL_ADDRESS_SIGNAL))) WHEN INSTRUCTION_COUNTER > 7;
	CONTROL_WORD(ROM_WIDTH-1 DOWNTO 23) <= ROM_OUTPUT(ROM_WIDTH-1 DOWNTO 23);
	CONTROL_WORD(14 DOWNTO 11) <= ROM_OUTPUT(14 DOWNTO 11);
	CONTROL_WORD(6 DOWNTO 0) <= ROM_OUTPUT(6 DOWNTO 0);
	-------------------------Place Holder circuits
	IR_SRC <= '0'&IR (8 DOWNTO 6);
	
	CONTROL_WORD(22 DOWNTO 19) <= STD_LOGIC_VECTOR(UNSIGNED (IR_SRC) + 1) WHEN ROM_OUTPUT(22 DOWNTO 19) = "1111"
		ELSE ROM_OUTPUT(22 DOWNTO 19) ;
	
	CONTROL_WORD(18 DOWNTO 15) <= STD_LOGIC_VECTOR(UNSIGNED (IR_SRC) + 1) WHEN ROM_OUTPUT(18 DOWNTO 15) = "1111"
		ELSE ROM_OUTPUT(18 DOWNTO 15) ;
	
	CONTROL_WORD(10 DOWNTO 7) <= STD_LOGIC_VECTOR(UNSIGNED (IR_SRC) + 1) WHEN ROM_OUTPUT(10 DOWNTO 7) = "1111"
		ELSE ROM_OUTPUT(10 DOWNTO 7) ;
	
END FETCH_SOURCE;
