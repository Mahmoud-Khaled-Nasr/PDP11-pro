LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE.ALL;

ENTITY IR_REGISTER IS
	GENERIC (SIZE : INTEGER := 16);
	PORT (
		CLK : IN STD_LOGIC;
		--THE SIZEOF THE IR IS 16 BIT ONLY
		DATA_IN : IN STD_LOGIC_VECTOR (SIZE-1 DOWNTO 0); 
		--USED TO ENABLE THE OUTPUT OF THE IR ON THE B BUS TO OUTPUT THE ADDRESS OF THE BRANCH
		BUS_B_OUT_ENABLE : IN STD_LOGIC ;
		BUS_B_IN_ENABLE : IN STD_LOGIC;
		DATA_OUT : OUT STD_LOGIC_VECTOR (SIZE+SIZE -1 DOWNTO 0)
	);
END ENTITY IR_REGISTER;
