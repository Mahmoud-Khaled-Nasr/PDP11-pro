LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE.ALL;

ENTITY IR_REGISTER IS
	GENERIC (IR_REG_SIZE : INTEGER := 32);
	PORT (
		D		: IN STD_LOGIC_VECTOR (IR_REG_SIZE-1 DOWNTO 0);	--DX : IF ENB=1 INPUT=D , IF ENBX=1 INPUT=DX
		CLK,RST,ENB	: IN STD_LOGIC;
		Q_BUS,Q_CU	: OUT STD_LOGIC_VECTOR (IR_REG_SIZE-1 DOWNTO 0)	--QX IS THE SAME AS 'Q' NO THING ELSE
	);

END ENTITY IR_REGISTER;


ARCHITECTURE IR_REGISTER_ARCH OF IR_REGISTER IS


BEGIN

process(RST,CLK,ENB)
	begin
		if (RST='1') then
			Q_bus<="00000000000000000000000000000001";
			Q_cu<="00000000000000000000000000000001";

		elsif(falling_edge(clk) and enb='1')then
			IF (D(7)='1') THEN
				Q_BUS <= "111111111111111111111111"&D(7 downto 0);
				Q_CU <= D;
			ELSE
				Q_BUS <= D;
				Q_CU <= D;
			END IF;
			
		end if;
	end process;


END IR_REGISTER_ARCH;