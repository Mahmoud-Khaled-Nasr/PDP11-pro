LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE.ALL;

ENTITY IR_REGISTER IS
	GENERIC (SIZE : INTEGER := 32);
	PORT (
		D		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);	--DX : IF ENB=1 INPUT=D , IF ENBX=1 INPUT=DX
		CLK,RST,ENB	: IN STD_LOGIC;
		Q 		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)	--QX IS THE SAME AS 'Q' NO THING ELSE
	);
END ENTITY IR_REGISTER;


ARCHITECTURE IR_REGISTER_ARCH OF IR_REGISTER IS


BEGIN

process(RST,CLK,ENB)
	begin
		if (RST='1') then
			Q<="00000000000000000000000000000001";
		elsif(falling_edge(clk) and enb='1')then
			Q<=D;
		end if;
	end process;


END IR_REGISTER_ARCH;