LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE;

ENTITY RAM IS
	GENERIC (ADDRESS_SIZE : INTEGER :=11; CELL_SIZE : INTEGER := 16*2);	--11BIT FOR MEMORY ADDRESS_SIZE PROVIDES 2K BIT MEMORY --16*2 : I ALLWAYS READ & WRITE 2 CELLS BUT I MAYBE WANT TO READ 1 CELL IN THIS CASE MDR WILL HANDLE IT
	PORT (
		DATA_IN 	:IN STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
		WRT	 	: IN STD_LOGIC;		
		CLK,ENB		:IN STD_LOGIC;					--RAM IS ALWAY ENABLED
		ADDRESS		:IN STD_LOGIC_VECTOR(ADDRESS_SIZE-1 DOWNTO 0);
		DATA_OUT 	: OUT STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
		--MDR_READ IS THE SIGNAL TO ENABLE THE MDR TO READ FROM THE MEMORY
		MFC, MDR_READ 	:OUT STD_LOGIC	--I DIDN'T USE THOSE SIGNALS TILL NOW
		
	);
END ENTITY RAM;
		

ARCHITECTURE RAM_ARCH OF RAM IS

	TYPE RAM_TYPE IS ARRAY(0 TO 2047) OF std_logic_vector(CELL_SIZE/2-1 DOWNTO 0);
	SIGNAL MEMORY : RAM_TYPE ;
	
	BEGIN
		PROCESS(CLK) IS
			BEGIN
				IF rising_edge(CLK) THEN  
					IF WRT = '1' THEN
						MEMORY(to_integer(unsigned(ADDRESS))) <= DATA_IN(15 DOWNTO 0);
						MEMORY(to_integer(unsigned(ADDRESS-1))) <= DATA_IN(CELL_SIZE-1 DOWNTO 16);
					END IF;
				END IF;
		END PROCESS;
		DATA_OUT(15 DOWNTO 0) <= MEMORY(to_integer(unsigned(ADDRESS)));
		DATA_OUT(CELL_SIZE-1 DOWNTO 16) <= MEMORY(to_integer(unsigned(ADDRESS-1)));

END RAM_ARCH;