LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE WORK.MY_PACKAGE.ALL;

ENTITY SRC_FETCHING_BLOCK IS
	--YOU CAN ADD ANY SIGNAL YOU WANT FOR EXAMPLE THE MODE OR OTHER SIGNALS
	PORT (
		IR : IN std_logic_vector (IR_SIZE-1 DOWNTO 0);
		INSTRUCTION_COUNTER : IN STD_LOGIC_VECTOR (INSTRUCTION_COUNTER_OUTPUT_SIZE-1 DOWNTO 0); 
		CONTROL_WORD: OUT STD_LOGIC_VECTOR (ROM_WIDTH-1 DOWNTO 0);
		INITIAL_ADDRESS: OUT STD_LOGIC_VECTOR (INSTRUCTION_COUNTER_OUTPUT_SIZE-1 DOWNTO 0) );
END ENTITY SRC_FETCHING_BLOCK;

ARCHITECTURE FETCH_SOURCE OF SRC_FETCHING_BLOCK IS
	
	-----------------ROM------------
	CONSTANT ROM_LENGTH : INTEGER := 5; --LENGTH OF THE ROM USED IN THIS BLOCK
	TYPE ROM_TYPE IS ARRAY(0 TO ROM_LENGTH - 1) OF std_logic_vector(ROM_WIDTH-1 DOWNTO 0);
	BEGIN
	-------------------------Circuit that calculate the initial value

	-------------------------the ROM process---------------

	-------------------------Other circuits
	--For example The Place holder cuircuit
	
	-- AT THE END ALL IS THE OUTPUT IS
	-- CONTROL_WORD <= SOMETHING RIGHT I HOPE
END FETCH_SOURCE;
